��/ /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     C o v e r a g e   C o l l e c t o r  
 / /   F i l e :         c o v e r a g e . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 6 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   S y s t e m V e r i l o g   c o v e r a g e   c o l l e c t o r   c l a s s   i s   r e s p o n s i b l e   f o r   g a t h e r i n g    
 / /   c o v e r a g e   i n f o r m a t i o n   f r o m   t h e   t r a n s a c t i o n s   i t   r e c e i v e s .  
 / /  
 / /   T h e   c o v e r a g e   c o l l e c t o r   c l a s s   h a s   a   t r a n s a c t i o n   o b j e c t   a n d   a   m a i l b o x    
 / /   ' d r i v 2 c o r ' ,   w h i c h   i s   u s e d   t o   r e c e i v e   t r a n s a c t i o n s   f r o m   t h e   d r i v e r .   I t   a l s o    
 / /   u s e s   a   v i r t u a l   i n t e r f a c e   ' v i f '   t o   c o m m u n i c a t e   w i t h   t h e   D U V .  
 / /  
 / /   T h e   c o v e r a g e   c o l l e c t o r   u s e s   a   c o v e r g r o u p   ' c o v _ c g '   t o   d e f i n e   t h e   c o v e r a g e    
 / /   p o i n t s   a n d   c r o s s e s   t h a t   i t   i s   i n t e r e s t e d   i n .   T h e   c o v e r a g e   p o i n t s   a r e    
 / /   t r a n s _ t y p e ,   H t r a n s ,   H s i z e ,   a n d   H b u r s t ,   w h i c h   a r e   p r o p e r t i e s   o f   t h e    
 / /   t r a n s a c t i o n .   T h e   c r o s s e s   a r e   c o m b i n a t i o n s   o f   t r a n s _ t y p e   w i t h   t h e   o t h e r    
 / /   p r o p e r t i e s .  
 / /  
 / /   T h e   ' e x e c u t e '   t a s k   i s   t h e   m a i n   r o u t i n e   o f   t h e   c o v e r a g e   c o l l e c t o r .   I t    
 / /   r e t r i e v e s   a   t r a n s a c t i o n   f r o m   t h e   d r i v e r   u s i n g   ' d r i v 2 c o r . g e t ( t x ) ' ,   a n d    
 / /   t h e n   i t   d i s p l a y s   i n f o r m a t i o n   a b o u t   t h e   t r a n s a c t i o n .  
 / /  
 / /   N o t e :   T h e   ' s a m p l e _ c o v e r a g e '   a n d   ' p r i n t _ c o v e r a g e '   f u n c t i o n s   a r e   c o m m e n t e d    
 / /   o u t   i n   t h e   o r i g i n a l   c o d e .   T h e   ' s a m p l e _ c o v e r a g e '   f u n c t i o n   w o u l d   b e   u s e d   t o    
 / /   s a m p l e   t h e   c o v e r a g e   p o i n t s   a n d   c r o s s e s   d e f i n e d   i n   ' c o v _ c g '   u s i n g   t h e   c u r r e n t    
 / /   t r a n s a c t i o n .   T h e   ' p r i n t _ c o v e r a g e '   f u n c t i o n   w o u l d   b e   u s e d   t o   p r i n t   a   c o v e r a g e    
 / /   r e p o r t ,   s h o w i n g   t h e   p e r c e n t a g e   o f   c o v e r a g e   p o i n t s   a n d   c r o s s e s   t h a t   h a v e   b e e n    
 / /   h i t .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
 c l a s s   c o v e r a g e _ c o l l e c t o r ;  
  
         T r a n s a c t i o n   t x ;           / /   T r a n s a c t i o n   o b j e c t  
         m a i l b o x   # ( T r a n s a c t i o n )   d r i v 2 c o r ;       / /   M a i l b o x   f o r   G e n e r a t o r   t o   D r i v e r  
         v i r t u a l   a h b _ a p b _ b f m _ i f   v i f ;  
         / /   C o v e r a g e   g r o u p s  
         c o v e r g r o u p   c o v _ c g ;  
                 t r a n s _ t y p e _ c p :   c o v e r p o i n t   t x . t r a n s _ t y p e   {  
                         b i n s   r e a d     =   { T r a n s a c t i o n : : A H B _ R E A D } ;  
                         b i n s   w r i t e   =   { T r a n s a c t i o n : : A H B _ W R I T E } ;  
                 }  
                 H t r a n s _ c p :   c o v e r p o i n t   t x . H t r a n s   {  
                         b i n s   n o n _ s e q   =   { 2 ' b 0 0 } ;  
                         b i n s   i d l e         =   { 2 ' b 0 1 } ;  
                         b i n s   s e q           =   { 2 ' b 1 0 } ;  
                         b i n s   b u s y         =   { 2 ' b 1 1 } ;  
                 }  
                 H s i z e _ c p :   c o v e r p o i n t   t x . H s i z e   {  
                         b i n s   s i z e _ b y t e           =   { 3 ' b 0 0 0 } ;  
                         b i n s   s i z e _ h a l f w o r d   =   { 3 ' b 0 0 1 } ;  
                         b i n s   s i z e _ w o r d           =   { 3 ' b 0 1 0 } ;  
                 }  
                 H b u r s t _ c p :   c o v e r p o i n t   t x . H b u r s t   {  
                         b i n s   s i n g l e   =   { 3 ' b 0 0 0 } ;  
                         b i n s   i n c r       =   { 3 ' b 0 0 1 } ;  
                         b i n s   w r a p 4     =   { 3 ' b 0 1 0 } ;  
                         b i n s   i n c r 4     =   { 3 ' b 0 1 1 } ;  
                 }  
                 / /   C r o s s   c o v e r a g e  
                 t r a n s _ x _ h t r a n s :   c r o s s   t r a n s _ t y p e _ c p ,   H t r a n s _ c p ;  
                 t r a n s _ x _ h s i z e :   c r o s s   t r a n s _ t y p e _ c p ,   H s i z e _ c p ;  
                 t r a n s _ x _ h b u r s t :   c r o s s   t r a n s _ t y p e _ c p ,   H b u r s t _ c p ;  
         e n d g r o u p  
  
         / /   c o v _ c g   a h b _ c g ;  
         f u n c t i o n   n e w ( m a i l b o x   # ( T r a n s a c t i o n )   d r i v 2 c o r ,   v i r t u a l   a h b _ a p b _ b f m _ i f   v i f ) ;  
                 t h i s . d r i v 2 c o r   =   d r i v 2 c o r ;  
               c o v _ c g   =   n e w ;  
                 t h i s . v i f   =   v i f ;  
         e n d f u n c t i o n  
  
         / /   F u n c t i o n   t o   s a m p l e   t h e   c o v e r a g e  
         / *   f u n c t i o n   v o i d   s a m p l e _ c o v e r a g e ( ) ;  
                 c o v _ c g . s a m p l e ( ) ;  
         e n d f u n c t i o n  
  
         / /   F u n c t i o n   t o   p r i n t   t h e   c o v e r a g e   r e p o r t  
         f u n c t i o n   v o i d   p r i n t _ c o v e r a g e ( ) ;  
                 $ d i s p l a y ( " C o v e r a g e :   % 0 d % % " ,   c o v _ c g . g e t _ c o v e r a g e ( )   *   1 0 0 ) ;  
         e n d f u n c t i o n   * /  
  
         / /   T a s k   t o   g e t   T r a n s a c t i o n   f r o m   m a i l b o x   a n d   s a m p l e   c o v e r a g e  
         t a s k   e x e c u t e ( ) ;  
                 f o r e v e r   b e g i n  
                         d r i v 2 c o r . g e t ( t x ) ;  
                       / /   s a m p l e _ c o v e r a g e ( ) ;  
                       $ d i s p l a y ( " t x   g o t " ,   t x ) ;  
                 e n d  
         e n d t a s k  
 e n d c l a s s  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     D r i v e r  
 / /   F i l e :         d r i v e r . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 6 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   S y s t e m V e r i l o g   d r i v e r   c l a s s   i s   r e s p o n s i b l e   f o r   r e c e i v i n g   t r a n s a c t i o n s    
 / /   f r o m   t h e   g e n e r a t o r   a n d   d r i v i n g   t h e m   i n t o   t h e   D e s i g n   U n d e r   V e r i f i c a t i o n   ( D U V ) .    
 / /   I t   c o m m u n i c a t e s   w i t h   t h e   D U V   t h r o u g h   a   v i r t u a l   i n t e r f a c e   ' v i f ' .  
 / /  
 / /   T h e   d r i v e r   c l a s s   h a s   t r a n s a c t i o n   h a n d l e s   a n d   s e v e r a l   m a i l b o x e s :   ' g e n 2 d r i v ' ,    
 / /   ' d r i v 2 s b ' ,   a n d   ' d r i v 2 c o r ' .   T h e   ' g e n 2 d r i v '   m a i l b o x   i s   u s e d   t o   r e c e i v e    
 / /   t r a n s a c t i o n s   f r o m   t h e   g e n e r a t o r ,   ' d r i v 2 s b '   s e n d s   t r a n s a c t i o n s   t o   t h e    
 / /   s c o r e b o a r d   f o r   v e r i f i c a t i o n ,   a n d   ' d r i v 2 c o r '   s e n d s   t r a n s a c t i o n s   d i r e c t l y    
 / /   t o   t h e   D U V .  
 / /  
 / /   T h e   ' d r i v e '   t a s k   i s   t h e   m a i n   r o u t i n e   o f   t h e   d r i v e r .   I t   r e t r i e v e s   a    
 / /   t r a n s a c t i o n   f r o m   t h e   g e n e r a t o r   u s i n g   ' g e n 2 d r i v . g e t ( t x ) ' ,   t h e n   s e n d s   i t    
 / /   t o   t h e   s c o r e b o a r d   a n d   t h e   D U V   u s i n g   ' d r i v 2 s b . p u t ( t x ) '   a n d   ' d r i v 2 c o r . p u t ( t x ) '    
 / /   r e s p e c t i v e l y .  
 / /  
 / /   A f t e r   t h a t ,   t h e   ' d r i v e '   t a s k   u s e s   t h e   v i r t u a l   i n t e r f a c e   t o   d r i v e   t h e    
 / /   t r a n s a c t i o n   v a l u e s   t o   t h e   D U V .   I t   a s s i g n s   e a c h   s i g n a l   i n   t h e   D U V   w i t h    
 / /   t h e   c o r r e s p o n d i n g   v a l u e   f r o m   t h e   t r a n s a c t i o n .   T h e n   i t   w a i t s   f o r   a   c l o c k    
 / /   e d g e   b e f o r e   p r o c e e d i n g .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
  
 c l a s s   d r i v e r ;  
  
         T r a n s a c t i o n   t x ;   / /   H a n d l e   f o r   t r a n s a c t i o n s                
  
         m a i l b o x   # ( T r a n s a c t i o n )   g e n 2 d r i v ;   / /   G e n e r a t o r   t o   D r i v e r   m a i l b o x  
         m a i l b o x   # ( T r a n s a c t i o n )   d r i v 2 s b ;     / /   D r i v e r   t o   S c o r e b o a r d   m a i l b o x  
         m a i l b o x   # ( T r a n s a c t i o n )   d r i v 2 c o r ;   / /   D r i v e r   t o   D U V   ( D e v i c e   U n d e r   V e r i f i c a t i o n )   m a i l b o x  
         v i r t u a l   a h b _ a p b _ b f m _ i f . m a s t e r   v i f ;                                   / /   V i r t u a l   i n t e r f a c e   t o   D U V  
  
         / /   C o n s t r u c t o r  
         f u n c t i o n   n e w ( m a i l b o x   # ( T r a n s a c t i o n ) g e n 2 d r i v ,   m a i l b o x   # ( T r a n s a c t i o n ) d r i v 2 s b ,   m a i l b o x   # ( T r a n s a c t i o n ) d r i v 2 c o r ,   v i r t u a l   a h b _ a p b _ b f m _ i f . m a s t e r   v i f ) ;  
                 t h i s . g e n 2 d r i v   =   g e n 2 d r i v ;   / /   a s s i g n i n g   g e n 2 d r i v    
                 t h i s . d r i v 2 s b   =   d r i v 2 s b ;       / /   a s s i g n i n g   d r i v 2 s b  
                 t h i s . d r i v 2 c o r   =   d r i v 2 c o r ;   / /   a s s i g n i n g   d r i v 2 c o r  
                 t h i s . v i f   =   v i f ;                       / /   a s s i g n i n g   v i r t u a l   i n t e r f a c e  
         e n d f u n c t i o n  
  
 / /   T a s k   t o   g e t   p a c k e t s   f r o m   g e n e r a t o r   a n d   d r i v e   t h e m   i n t o   i n t e r f a c e  
 t a s k   d r i v e ;    
         g e n 2 d r i v . g e t ( t x ) ;        
         d r i v 2 s b . p u t ( t x ) ;        
         d r i v 2 c o r . p u t ( t x ) ;  
         $ d i s p l a y ( " d r i v e r   t x " ,   t x ) ;  
         / /   D r i v i n g   t h e   v a l u e s   t o   t h e   D U V   v i a   t h e   v i r t u a l   i n t e r f a c e  
         v i f . d r v _ c b . H w r i t e   < =   t x . H w r i t e ;            
         v i f . d r v _ c b . H t r a n s   < =   t x . H t r a n s ;  
         v i f . d r v _ c b . H w d a t a   < =   t x . H w d a t a ;            
         v i f . d r v _ c b . H a d d r   < =   t x . H a d d r ;  
       # 1 0 ;     / /   w a i t   f o r   1 0   t i m e   u n i t s  
         / /   v i f . d r v _ c b . H s i z e   < =   t x . H s i z e ;              
         / /   v i f . d r v _ c b . H b u r s t   < =   t x . H b u r s t ;          
 e n d t a s k  
 e n d c l a s s  
  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     E n v i r o n m e n t  
 / /   F i l e :         e n v i r o n m e n t . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 9 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   e n v i r o n m e n t   c l a s s   i s   a   c e n t r a l   p a r t   o f   t h e   v e r i f i c a t i o n   p r o c e s s   i n   a    
 / /   S y s t e m V e r i l o g   t e s t b e n c h .   I t   h o u s e s   a l l   t h e   m a i n   v e r i f i c a t i o n   c o m p o n e n t s   s u c h    
 / /   a s   t h e   g e n e r a t o r ,   d r i v e r ,   m o n i t o r ,   a n d   s c o r e b o a r d ,   a n d   m a n a g e s   t h e   i n t e r a c t i o n s    
 / /   b e t w e e n   t h e m .    
 / /   I n   t h i s   p a r t i c u l a r   s c e n a r i o ,   i t   e s t a b l i s h e s   m a i l b o x e s   f o r   c o m m u n i c a t i o n ,    
 / /   i n i t i a t e s   a l l   c o m p o n e n t s ,   a n d   m a n a g e s   s p e c i f i c   t e s t   c a s e s .   T h e s e   t e s t   c a s e s    
 / /   r e p r e s e n t   v a r i o u s   t r a n s a c t i o n s   t h a t   t h e   A H B   A P B   b r i d g e   s h o u l d   b e   c a p a b l e   o f    
 / /   h a n d l i n g ,   t h u s   f a c i l i t a t i n g   c o m p r e h e n s i v e   t e s t i n g   a n d   v e r i f i c a t i o n   o f   t h e    
 / /   d e s i g n   u n d e r   t e s t   ( D U T ) .  
 / /  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
  
 c l a s s   e n v i r o n m e n t ;  
     m a i l b o x   # ( T r a n s a c t i o n )   g e n 2 d r i v ;      
     m a i l b o x   # ( T r a n s a c t i o n )   d r i v 2 s b ;      
     m a i l b o x   # ( T r a n s a c t i o n )   m a i l 2 s b ;    
     m a i l b o x   # ( T r a n s a c t i o n )   d r i v 2 c o r ;  
  
     g e n e r a t o r   g e n ;                  
     d r i v e r   d r i v ;                      
     a h b _ a p b _ m o n i t o r   m o n i ;                    
     a h b _ a p b _ s c o r e b o a r d   s b ;                  
     / /   c o v e r a g e _ c o l l e c t o r   c o v ;  
     v i r t u a l   a h b _ a p b _ b f m _ i f   v i f ;  
  
     f u n c t i o n   n e w ( v i r t u a l   a h b _ a p b _ b f m _ i f   v i f ) ;  
         t h i s . v i f   =   v i f ;  
     e n d f u n c t i o n  
  
     f u n c t i o n   c r e a t e ( ) ;  
         g e n 2 d r i v   =   n e w ( 1 ) ;  
         d r i v 2 s b   =   n e w ( 1 ) ;  
         m a i l 2 s b   =   n e w ( 1 ) ;  
         d r i v 2 c o r   =   n e w ( 1 ) ;  
         g e n   =   n e w ( g e n 2 d r i v ) ;  
         d r i v   =   n e w ( g e n 2 d r i v ,   d r i v 2 s b ,   d r i v 2 c o r ,   v i f ) ;  
         m o n i   =   n e w ( m a i l 2 s b ,   v i f ) ;  
         s b   =   n e w ( d r i v 2 s b ,   m a i l 2 s b ) ;  
         / /   c o v   =   n e w ( d r i v 2 c o r ,   v i f ) ;  
     e n d f u n c t i o n  
  
 / *  
     t a s k   e n v _ r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
         f o r k  
             g e n . w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
             d r i v . d r i v e ( ) ;  
             m o n i . w a t c h ( ) ;  
             s b . d a t a _ w r i t e ( ) ;  
  
         j o i n _ n o n e  
     e n d t a s k  
  
 * /  
  
 	 / /   T e s t   C a s e   2  
 t a s k   e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3  
 t a s k   e n v _ r e a d _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4  
 t a s k   e n v _ w r i t e _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5  
 t a s k   e n v _ r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   6  
 t a s k   e n v _ w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   7  
 t a s k   e n v _ r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   8  
 t a s k   e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   9  
 t a s k   e n v _ r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 0  
 t a s k   e n v _ w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 1  
 t a s k   e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 2  
 t a s k   e n v _ w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 3  
 t a s k   e n v _ r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 4  
 t a s k   e n v _ w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 5  
 t a s k   e n v _ r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 6  
 t a s k   e n v _ w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
 $ d i s p l a y ( " i n   e n v " ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 7  
 t a s k   e n v _ r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 8  
 t a s k   e n v _ w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   1 9  
 t a s k   e n v _ r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 0  
 t a s k   e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 1  
 t a s k   e n v _ r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 2  
 t a s k   e n v _ w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 3  
 t a s k   e n v _ r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 4  
 t a s k   e n v _ w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 5  
 t a s k   e n v _ r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 6  
 t a s k   e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 7  
 t a s k   e n v _ r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 8  
 t a s k   e n v _ w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   2 9  
 t a s k   e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 0  
 t a s k   e n v _ w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 1  
 t a s k   e n v _ r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 2  
 t a s k   e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 3  
 t a s k   e n v _ r e a d _ s i n g l e _ w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / / h e r e  
 / /   T e s t   C a s e   3 4  
 t a s k   e n v _ w r i t e _ i n c r _ b y t e _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r _ b y t e _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 5  
 t a s k   e n v _ r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 6  
 t a s k   e n v _ w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 7  
 t a s k   e n v _ r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 8  
 t a s k   e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   3 9  
 t a s k   e n v _ r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 0  
 t a s k   e n v _ w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 1  
 t a s k   e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 2  
 t a s k   e n v _ w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 3  
 t a s k   e n v _ r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 4  
 t a s k   e n v _ w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 5  
 t a s k   e n v _ r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 6  
 t a s k   e n v _ w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 7  
 t a s k   e n v _ r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 8  
 t a s k   e n v _ w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   4 9  
 t a s k   e n v _ r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 0  
 t a s k   e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 1  
 t a s k   e n v _ r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 2  
 t a s k   e n v _ w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 3  
 t a s k   e n v _ r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 4  
 t a s k   e n v _ w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 5  
 t a s k   e n v _ r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 6  
 t a s k   e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 7  
 t a s k   e n v _ r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 8  
 t a s k   e n v _ w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   5 9  
 t a s k   e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ r e a d ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   6 0  
 t a s k   e n v _ w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   6 1  
 t a s k   e n v _ w r i t e _ i n c r 4 _ w o r d _ i d l e _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ w o r d _ i d l e _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   6 2  
 t a s k   e n v _ w r i t e _ i n c r 4 _ w o r d _ b u s y _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
     f o r k  
         g e n . w r i t e _ i n c r 4 _ w o r d _ b u s y _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 / /   T e s t   C a s e   6 3  
 t a s k   e n v _ w r i t e _ s i n g l e _ b y t e _ i d l e _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
     f o r k  
         g e n . w r i t e _ s i n g l e _ b y t e _ i d l e _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
         d r i v . d r i v e ( ) ;  
         m o n i . w a t c h ( ) ;  
         s b . d a t a _ w r i t e ( ) ;  
     j o i n _ n o n e  
 e n d t a s k  
  
 e n d c l a s s  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     G e n e r a t o r  
 / /   F i l e :         g e n e r a t o r . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 9 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   S y s t e m V e r i l o g   g e n e r a t o r   c l a s s   g e n e r a t e s   t r a n s a c t i o n s   o f   d i f f e r e n t    
 / /   t y p e s   a n d   s e n d s   t h e m   t o   t h e   d r i v e r   f o r   e x e c u t i o n .   I n   t h i s   m o d u l e ,   t h e r e    
 / /   a r e   s e v e r a l   t e s t   c a s e s   d e f i n e d   a s   t a s k s ,   e a c h   r e p r e s e n t i n g   a   u n i q u e    
 / /   t r a n s a c t i o n .  
 / /  
 / /   T h e   c l a s s   g e n e r a t o r   h a s   a   t r a n s a c t i o n   h a n d l e   ' t x '   a n d   a   m a i l b o x   ' g e n 2 d r i v '  
 / /   t h a t   i s   u s e d   t o   s e n d   t r a n s a c t i o n s   t o   t h e   d r i v e r .   I t   a l s o   h a s   a   v i r t u a l  
 / /   i n t e r f a c e   ' v i f '   t o   c o m m u n i c a t e   w i t h   t h e   D U T .  
 / /  
 / /   T h e   ' r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y '   t a s k ,   f o r   i n s t a n c e ,    
 / /   c r e a t e s   a   r e a d   t r a n s a c t i o n ,   w i t h   e a c h   f i e l d   o f   t h e   t r a n s a c t i o n   b e i n g    
 / /   a s s i g n e d   a   v a l u e   a c c o r d i n g   t o   t h e   r e q u i r e m e n t s   o f   t h e   t e s t   c a s e .   O n c e   t h e    
 / /   t r a n s a c t i o n   i s   r e a d y ,   i t   i s   s e n t   t o   t h e   d r i v e r   u s i n g   t h e   ' g e n 2 d r i v . p u t ( t x ) ; '    
 / /   c o m m a n d .  
 / /  
 / /   S i m i l a r   o p e r a t i o n s   a r e   p e r f o r m e d   i n   o t h e r   t e s t   c a s e   t a s k s .   E a c h   t a s k    
 / /   d e f i n e s   a   d i f f e r e n t   t y p e   o f   t r a n s a c t i o n ,   w i t h   v a r i o u s   v a l u e s   a s s i g n e d   t o    
 / /   t h e   f i e l d s   o f   t h e   t r a n s a c t i o n .  
 / /  
 / /   T h e   g e n e r a t o r   c l a s s   a l s o   s a m p l e s   e a c h   t r a n s a c t i o n   f o r   c o v e r a g e   u s i n g   t h e    
 / /   ' t x . c o v _ c g . s a m p l e ( ) ; '   c o m m a n d .   T h i s   h e l p s   t o   e n s u r e   t h a t   a l l   t y p e s   o f    
 / /   t r a n s a c t i o n s   a r e   g e n e r a t e d   a n d   e x e c u t e d ,   t h u s   e n s u r i n g   c o m p l e t e   f u n c t i o n a l    
 / /   c o v e r a g e .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
 c l a s s   g e n e r a t o r ;  
  
         T r a n s a c t i o n   t x ;       / /   H a n d l e   f o r   H t r a n s a c t i o n s                      
         m a i l b o x   # ( T r a n s a c t i o n )   g e n 2 d r i v ;     / /   G e n e r a t o r   t o   D r i v e r   m a i l b o x  
  
         l o g i c   [ 3 1 : 0 ]   t e m p _ H a d d r ;   / /   t e m p o r a r y   v a r i a b l e      
         l o g i c   [ 1 1 : 0 ]   H a d d r _ a r r a y   [ 6 ]   =     { 8 ' h 1 1 ,   8 ' h 2 2 ,   1 2 ' h 3 8 4 ,   1 2 ' h F D 2 ,   1 2 ' h 6 4 ,   1 2 ' h D A C } ;   / /   H a d d r e s s   a r r a y  
         l o g i c   [ 1 1 : 0 ]   H a d d r _ H b u r s t [ 2 ]   =   { 1 2 ' h a b   ,   1 2 ' h d e } ;   / /   H b u r s t  
         i n t   i   = 0 ;  
  
         f u n c t i o n   n e w ( m a i l b o x   # ( T r a n s a c t i o n ) g e n 2 d r i v ) ;  
                 t h i s . g e n 2 d r i v       =   g e n 2 d r i v ;  
         e n d f u n c t i o n  
          
         / /   T e s t   C a s e   2  
         t a s k   w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;   / /   W r i t e   o p e r a t i o n  
         t x . u p d a t e _ t r a n s _ t y p e ( ) ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
         t x . P e n a b l e   =   1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;   / /   G e n e r a t e   r a n d o m   d a t a   f o r   w r i t e  
         t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
  
         / /   T e s t   C a s e   3  
         t a s k   r e a d _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
         t x . P e n a b l e   =   1 ;  
         t x . P w r i t e   =   0 ;  
         t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
             t x . u p d a t e _ t r a n s _ t y p e ( ) ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4  
         t a s k   w r i t e _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ e r r o r   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s p   =   1 ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
     	 t x . u p d a t e _ t r a n s _ t y p e ( ) ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5  
         t a s k   r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   6  
         t a s k   w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . P e n a b l e   =   1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   7  
         t a s k   r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   8  
         t a s k   w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   9  
         t a s k   r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 0  
         t a s k   w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 1  
         t a s k   r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . P e n a b l e   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 2  
         t a s k   w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 3  
         t a s k   r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 4  
         t a s k   w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 1 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 5  
         t a s k   r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 6  
         t a s k   w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 7  
         t a s k   r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 1 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 8  
         t a s k   w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   1 9  
         t a s k   r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 0  
         t a s k   w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 1  
         t a s k   r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 2  
         t a s k   w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s p   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 3  
         t a s k   r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 4  
         t a s k   w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 5  
         t a s k   r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 6  
         t a s k   w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 7  
         t a s k   r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 8  
         t a s k   w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   2 9  
         t a s k   r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 0  
         t a s k   w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 1  
         t a s k   r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 2  
         t a s k   w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 3  
         t a s k   r e a d _ s i n g l e _ w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 4  
         t a s k   w r i t e _ i n c r _ b y t e _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r _ b y t e _ n o n s e q _ i n c r _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 5  
         t a s k   r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 6  
         t a s k   w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 7  
         t a s k   r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 8  
         t a s k   w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   3 9  
         t a s k   r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 0  
         t a s k   w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 1  
         t a s k   r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 2  
         t a s k   w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 3  
         t a s k   r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 4  
         t a s k   w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
     	 t x . t r a n s _ t y p e   =   T r a n s a c t i o n : : A H B _ W R I T E ;   / /   S e t   t r a n s a c t i o n   t y p e   a s   W R I T E  
  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 1 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 5  
         t a s k   r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 6  
         t a s k   w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 7  
         t a s k   r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 1 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 8  
         t a s k   w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 1 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   4 9  
         t a s k   r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 0  
         t a s k   w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 1  
         t a s k   r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 2  
         t a s k   w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s p   =   1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 3  
         t a s k   r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 4  
         t a s k   w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 5  
         t a s k   r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 6  
         t a s k   w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 7  
         t a s k   r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 0 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 8  
         t a s k   w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   5 9  
         t a s k   r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   0 ;  
                 t x . H s i z e   =   3 ' b 0 0 1 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   6 0  
         t a s k   w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 1 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   6 1  
         t a s k   w r i t e _ i n c r 4 _ w o r d _ i d l e _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ w o r d _ i d l e _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 0 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   6 2  
         t a s k   w r i t e _ i n c r 4 _ w o r d _ b u s y _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ i n c r 4 _ w o r d _ b u s y _ i n c r 4 _ H b u r s t _ r e s e t   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 1 0 ;  
                 t x . H b u r s t   =   3 ' b 0 1 1 ;  
                 t x . H t r a n s   =   2 ' b 0 1 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s e t   =   1 ;  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
         / /   T e s t   C a s e   6 3  
         t a s k   w r i t e _ s i n g l e _ b y t e _ i d l e _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
                 $ d i s p l a y ( $ t i m e ,   "       w r i t e _ s i n g l e _ b y t e _ i d l e _ s i n g l e _ H t r a n s f e r _ e r r o r   t a s k   i n   g e n e r a t o r " ) ;  
                 t x   =   n e w ( ) ;  
                 t x . H a d d r   =   $ u r a n d o m ;  
                 t x . H w r i t e   =   1 ;  
                 t x . H s i z e   =   3 ' b 0 0 0 ;  
                 t x . H b u r s t   =   3 ' b 0 0 0 ;  
                 t x . H t r a n s   =   2 ' b 0 0 ;  
                 t x . H w d a t a   =   $ u r a n d o m ( ) ;  
                 t x . h r e s p   =   1 ;  
 	 t x . c o v _ c g . s a m p l e ( ) ;   / /   A f t e r   t r a n s a c t i o n   i s   f u l l y   d e f i n e d  
                 g e n 2 d r i v . p u t ( t x ) ;  
         e n d t a s k  
  
 e n d c l a s s  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     I n t e r f a c e  
 / /   F i l e :         i n t e r f a c e . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 5 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   S y s t e m V e r i l o g   i n t e r f a c e   e n c a p s u l a t e s   t h e   s i g n a l s   o f   a   s p e c i f i c   p r o t o c o l    
 / /   ( i n   t h i s   c a s e   A H B - A P B   B r i d g e   p r o t o c o l )   a n d   p r o v i d e s   a   s i n g l e   h a n d l e   t o    
 / /   m a n a g e   t h e s e   s i g n a l s .   I t   a l s o   h e l p s   i n   e s t a b l i s h i n g   c o m m u n i c a t i o n   b e t w e e n    
 / /   d i f f e r e n t   v e r i f i c a t i o n   c o m p o n e n t s ,   l i k e   d r i v e r ,   m o n i t o r ,   a n d   D U T .  
 / /  
 / /   I n   t h i s   m o d u l e ,   t h e r e   a r e   t w o   c l o c k i n g   b l o c k s   d e f i n e d   f o r   t h e   d r i v e r   a n d    
 / /   m o n i t o r .   C l o c k i n g   b l o c k s   a l l o w   p r e c i s e   c o n t r o l   o v e r   w h e n   s i g n a l s   a r e   d r i v e n    
 / /   o r   s a m p l e d ,   w h i c h   i s   c r u c i a l   i n   d e s i g n   a n d   v e r i f i c a t i o n .  
 / /  
 / /   T h e   ' d r v _ c b '   b l o c k   i s   u s e d   b y   t h e   d r i v e r   t o   d r i v e   s i g n a l s   t o   t h e   D U T .   O n   t h e    
 / /   o t h e r   h a n d ,   t h e   ' m o n _ c b '   b l o c k   i s   u s e d   b y   t h e   m o n i t o r   t o   s a m p l e   s i g n a l s   f r o m    
 / /   t h e   D U T .   T h i s   w a y ,   w e   e n s u r e   t h a t   b o t h   t h e   d r i v e r   a n d   m o n i t o r   a r e   o p e r a t i n g    
 / /   s y n c h r o n o u s l y   w i t h   t h e   c l o c k .  
 / /  
 / /   T h e   m o d p o r t s   ' m a s t e r '   a n d   ' s l a v e '   a r e   d e f i n e d   t o   r e p r e s e n t   t h e   v i e w s   o f   t h e    
 / /   d r i v e r   a n d   m o n i t o r ,   r e s p e c t i v e l y .   T h e   d r i v e r   ( m a s t e r )   d r i v e s   t h e   s i g n a l s ,    
 / /   w h e r e a s   t h e   m o n i t o r   ( s l a v e )   s a m p l e s   t h e   s i g n a l s .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
  
 i n t e r f a c e   a h b _ a p b _ b f m _ i f ( i n p u t   w i r e   c l k ,   r e s e t n ) ;  
  
     / /   A H B   s i g n a l s  
     l o g i c   H w r i t e ;           / /   A H B   w r i t e   s i g n a l  
     l o g i c   H r e a d y i n ;       / /   A H B   r e a d y   i n p u t   s i g n a l  
     l o g i c   [ 1 : 0 ]   H t r a n s ;   / /   A H B   t r a n s f e r   t y p e   e n c o d i n g  
     l o g i c   [ 3 1 : 0 ]   H w d a t a ;   / /   A H B   w r i t e   d a t a  
     l o g i c   [ 3 1 : 0 ]   H a d d r ;     / /   A H B   a d d r e s s  
     l o g i c   [ 3 1 : 0 ]   H r d a t a ;   / /   A H B   r e a d   d a t a  
     l o g i c   [ 1 : 0 ]   H r e s p ;       / /   A H B   r e s p o n s e  
     l o g i c   H r e a d y o u t ;           / /   A H B   r e a d y   o u t p u t   s i g n a l  
  
     / /   A P B   s i g n a l s  
     w i r e   P e n a b l e ;               / /   A P B   e n a b l e   s i g n a l  
     w i r e   P w r i t e ;                 / /   A P B   w r i t e   s i g n a l  
     w i r e   [ 2 : 0 ]   P s e l x ;       / /   A P B   s e l e c t   s i g n a l s  
     w i r e   [ 3 1 : 0 ]   P w d a t a ;   / /   A P B   w r i t e   d a t a  
     w i r e   [ 3 1 : 0 ]   P a d d r ;     / /   A P B   a d d r e s s  
     w i r e   [ 3 1 : 0 ]   P r d a t a ;   / /   A P B   r e a d   d a t a  
  
     / /   C l o c k i n g   b l o c k   f o r   d r i v e r  
     / /   T h i s   b l o c k   d e f i n e s   t h e   t i m i n g   o f   t h e   s i g n a l s   w h e n   t h e y   a r e   d r i v e n   b y   t h e   d r i v e r  
     c l o c k i n g   d r v _ c b   @ ( p o s e d g e   c l k ) ;  
         d e f a u l t   i n p u t   # 1 n s   o u t p u t   # 1 n s ;   / /   D e f a u l t   s k e w   f o r   i n p u t   a n d   o u t p u t   s i g n a l s  
         o u t p u t   H w r i t e ,   H r e a d y i n ,   H t r a n s ,   H w d a t a ,   H a d d r ;   / /   A H B   s i g n a l s   d r i v e n   b y   t h e   d r i v e r  
         o u t p u t   P e n a b l e ,   P w r i t e ,   P s e l x ,   P w d a t a ,   P a d d r ;       / /   A P B   s i g n a l s   d r i v e n   b y   t h e   d r i v e r  
     e n d c l o c k i n g  
  
     / /   C l o c k i n g   b l o c k   f o r   m o n i t o r  
     / /   T h i s   b l o c k   d e f i n e s   t h e   t i m i n g   o f   t h e   s i g n a l s   w h e n   t h e y   a r e   m o n i t o r e d  
     c l o c k i n g   m o n _ c b   @ ( p o s e d g e   c l k ) ;  
         d e f a u l t   i n p u t   # 1 n s   o u t p u t   # 1 n s ;   / /   D e f a u l t   s k e w   f o r   i n p u t   a n d   o u t p u t   s i g n a l s  
         i n p u t   H w r i t e ,   H r e a d y i n ,   H t r a n s ,   H w d a t a ,   H a d d r ,   H r d a t a ,   H r e s p ,   H r e a d y o u t ;   / /   A H B   s i g n a l s   m o n i t o r e d  
         i n p u t   P e n a b l e ,   P w r i t e ,   P s e l x ,   P w d a t a ,   P a d d r ,   P r d a t a ;   / /   A P B   s i g n a l s   m o n i t o r e d  
     e n d c l o c k i n g  
  
     / /   M o d p o r t s  
     / /   T h e s e   d e f i n e   t h e   i n t e r f a c e   f o r   t h e   d r i v e r   a n d   m o n i t o r ,   r e s p e c t i v e l y  
     m o d p o r t   m a s t e r ( c l o c k i n g   d r v _ c b ,   i n p u t   c l k ,   r e s e t n ) ;   / /   d r i v e r  
     m o d p o r t   s l a v e ( c l o c k i n g   m o n _ c b ,   i n p u t   c l k ,   r e s e t n ) ;   / /   m o n i t o r  
  
 e n d i n t e r f a c e  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     M o n i t o r  
 / /   F i l e :         m o n i t o r . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 9 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   m o n i t o r   c l a s s   i s   a   c r u c i a l   p a r t   o f   t h e   v e r i f i c a t i o n   p r o c e s s   i n   a    
 / /   S y s t e m V e r i l o g   t e s t b e n c h .   I t   o b s e r v e s   t h e   i n t e r f a c e ,   c a p t u r e s   t h e    
 / /   t r a n s a c t i o n s   o c c u r r i n g   o n   t h e   b u s ,   a n d   f o r w a r d s   t h e m   t o   t h e   s c o r e b o a r d   f o r    
 / /   c h e c k i n g   a g a i n s t   t h e   e x p e c t e d   r e s u l t s .   I t   a c t s   a s   a   l i s t e n e r ,   m a k i n g   i t    
 / /   p a s s i v e   a n d   n o n - i n t r u s i v e   t o   t h e   d e s i g n   u n d e r   t e s t   ( D U T ) .  
 / /  
 / /   I n   t h i s   p a r t i c u l a r   s c e n a r i o ,   t h e   m o n i t o r   w a t c h e s   t h e   s i g n a l s   o n   t h e   A H B   A P B    
 / /   b r i d g e   i n t e r f a c e ,   c r e a t e s   t r a n s a c t i o n   o b j e c t s   r e p r e s e n t i n g   t h e   o b s e r v e d    
 / /   t r a n s a c t i o n s ,   a n d   s e n d s   t h e m   t o   t h e   s c o r e b o a r d .   I t   o p e r a t e s   i n   a n   i n f i n i t e    
 / /   l o o p ,   c o n t i n u o u s l y   m o n i t o r i n g   t h e   i n t e r f a c e   f o r   n e w   t r a n s a c t i o n s .  
 / /  
 / /   T h e   m o n i t o r   u t i l i z e s   a   c l o c k i n g   b l o c k   ( m o n _ c b )   t o   s a m p l e   t h e   i n t e r f a c e    
 / /   s i g n a l s   s y n c h r o n o u s l y   w i t h   t h e   c l o c k .   T h e   s a m p l e d   v a l u e s   a r e   u s e d   t o   c r e a t e    
 / /   t h e   t r a n s a c t i o n   o b j e c t ,   w h i c h   i s   t h e n   f o r w a r d e d   t o   t h e   s c o r e b o a r d   v i a   a    
 / /   m a i l b o x .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
 c l a s s   a h b _ a p b _ m o n i t o r ;  
  
         T r a n s a c t i o n   t x ;             / /   T r a n s a c t i o n   h a n d l e                          
         m a i l b o x   # ( T r a n s a c t i o n )   m a i l 2 s b ;     / /   M a i l b o x   t o   t h e   s c o r e b o a r d  
  
         / /   V i r t u a l   i n t e r f a c e   r e f e r e n c e  
         v i r t u a l   a h b _ a p b _ b f m _ i f . s l a v e   v i f ;                          
          
         f u n c t i o n   n e w ( m a i l b o x   # ( T r a n s a c t i o n )   m a i l 2 s b ,   v i r t u a l   a h b _ a p b _ b f m _ i f . s l a v e   v i f ) ;  
                 t h i s . m a i l 2 s b   =   m a i l 2 s b ;  
                 t h i s . v i f   =   v i f ;  
         e n d f u n c t i o n  
  
         / /   W a t c h   a n d   s e n d   t r a n s a c t i o n s   t o   t h e   s c o r e b o a r d  
         t a s k   w a t c h ;  
                 t x   =   n e w ( ) ;  
                  
                 / /   L o o p   t o   m o n i t o r   t r a n s a c t i o n s  
                 f o r e v e r   b e g i n  
                         @ ( v i f . m o n _ c b )   b e g i n     / /   U s e   t h e   c l o c k i n g   b l o c k   t o   s a m p l e   t h e   i n t e r f a c e   s i g n a l s  
                                 w a i t ( v i f . m o n _ c b . H t r a n s   ! = =   2 ' b 0 0 ) ;   / /   W a i t   f o r   a n y   t r a n s a c t i o n   t o   s t a r t  
                                 / / t x . t r a n s _ t y p e   =   v i f . m o n _ c b . H w r i t e   ?   T r a n s a c t i o n . A H B _ W R I T E   :   T r a n s a c t i o n . A H B _ R E A D ;  
                                 t x . H a d d r             =   v i f . m o n _ c b . H a d d r ;  
                                 t x . H w d a t a           =   v i f . m o n _ c b . H w d a t a ;  
                                 t x . H w r i t e           =   v i f . m o n _ c b . H w r i t e ;  
                                 t x . H t r a n s           =   v i f . m o n _ c b . H t r a n s ;  
                                 t x . P a d d r             =   v i f . m o n _ c b . P a d d r ;  
                                 t x . P w d a t a           =   v i f . m o n _ c b . P w d a t a ;  
                                 t x . P w r i t e           =   v i f . m o n _ c b . P w r i t e ;  
                                 t x . P s e l x             =   v i f . m o n _ c b . P s e l x ;  
                                 t x . P r d a t a           =   v i f . m o n _ c b . P r d a t a ;  
                                  
                                 m a i l 2 s b . p u t ( t x ) ;   / /   S e n d   t h e   t r a n s a c t i o n   t o   t h e   s c o r e b o a r d  
                         e n d  
                 e n d  
         e n d t a s k  
  
 e n d c l a s s  
  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     S c o r e b o a r d  
 / /   F i l e :         s c o r e b o a r d . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 6 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   S c o r e b o a r d   c l a s s   p l a y s   a   c r u c i a l   r o l e   i n   v e r i f i c a t i o n   p r o c e s s   a s   i t    
 / /   v a l i d a t e s   t h e   c o r r e c t n e s s   o f   t h e   d e s i g n .   I t   c o n t a i n s   a   m e m o r y   m o d e l   t h a t  
 / /   m i m i c s   t h e   b e h a v i o u r   o f   t h e   d e s i g n   u n d e r   t e s t   ( D U T ) .  
 / /  
 / /   T h e   S c o r e b o a r d   r e c e i v e s   t r a n s a c t i o n s   f r o m   b o t h   t h e   d r i v e r   a n d   t h e   m o n i t o r ,    
 / /   a l l o w i n g   i t   t o   c o m p a r e   t h e   e x p e c t e d   a n d   a c t u a l   r e s p o n s e s .   T h i s   c l a s s   h a s    
 / /   m e t h o d s   t o   h a n d l e   b o t h   d a t a   w r i t e   a n d   r e a d   o p e r a t i o n s .   F o r   a   w r i t e   o p e r a t i o n ,    
 / /   i t   v e r i f i e s   t h a t   t h e   d a t a   h a s   b e e n   c o r r e c t l y   w r i t t e n   i n t o   t h e   m e m o r y   m o d e l .    
 / /   F o r   a   r e a d   o p e r a t i o n ,   i t   c h e c k s   i f   t h e   d a t a   r e a d   f r o m   t h e   D U T   m a t c h e s   w i t h    
 / /   t h e   d a t a   s t o r e d   i n   t h e   m e m o r y   m o d e l .   A n y   d i s c r e p a n c y   i n   d a t a   w o u l d   r e s u l t    
 / /   i n   a n   a s s e r t i o n   e r r o r ,   f l a g g i n g   a   f a i l u r e   i n   t h e   v e r i f i c a t i o n   p r o c e s s .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
 c l a s s   a h b _ a p b _ s c o r e b o a r d ;  
  
         T r a n s a c t i o n   t x 1 ,   t x 2 ;  
         m a i l b o x   # ( T r a n s a c t i o n )   d r v 2 s b ;  
         m a i l b o x   # ( T r a n s a c t i o n )   m a i l 2 s b ;  
         l o g i c   [ 1 9 : 0 ]   t e m p _ a d d r ;   / /   W e   w i l l   o n l y   t r a c k   t h e   l e a s t   s i g n i f i c a n t   2 0   b i t s  
  
         b i t   [ 3 1 : 0 ]   m e m _ t b   [ 2 * * 2 0 ] ;   / /   m e m o r y   o f   2 ^ 2 0   l o c a t i o n s   e a c h   o f   3 2   b i t s  
  
         f u n c t i o n   n e w ( m a i l b o x   # ( T r a n s a c t i o n )   d r v 2 s b ,   m a i l b o x   # ( T r a n s a c t i o n )   m a i l 2 s b ) ;  
                 t h i s . d r v 2 s b   =   d r v 2 s b ;  
                 t h i s . m a i l 2 s b   =   m a i l 2 s b ;  
         e n d f u n c t i o n  
  
         t a s k   d a t a _ w r i t e ( ) ;  
  
                 $ d i s p l a y ( " S c o r e b o a r d   c h e c k . . . " ) ;  
  
                 / /   R e c e i v e   d a t a   f r o m   d r i v e r   a n d   m o n i t o r  
                 d r v 2 s b . g e t ( t x 1 ) ;  
                 m a i l 2 s b . g e t ( t x 2 ) ;  
  
                 t e m p _ a d d r   =   t x 1 . H a d d r [ 1 9 : 0 ] ;  
  
                 / /   W r i t e   d a t a   t o   t h e   m e m o r y   m o d e l  
                 m e m _ t b [ t e m p _ a d d r ]   =   t x 1 . H w d a t a ;  
  
                 $ d i s p l a y ( " I n p u t   A d d r e s s :   % h " ,   t e m p _ a d d r ) ;  
                 $ d i s p l a y ( " I n p u t   W r i t e   D a t a :   % h " ,   t x 1 . H w d a t a ) ;  
                 $ d i s p l a y ( " D a t a   S t o r e d :   % h " ,   m e m _ t b [ t e m p _ a d d r ] ) ;  
  
                 / /   A s s e r t   t h a t   t h e   d a t a   w a s   w r i t t e n   c o r r e c t l y  
                         a s s e r t   ( t x 1 . H w d a t a   = =   m e m _ t b [ t e m p _ a d d r ] )  
                         e l s e   $ e r r o r ( " D a t a   f a i l e d   t o   w r i t e " ) ;  
  
                 $ d i s p l a y ( " " ) ;  
 	 # 1 0 ;  
         e n d t a s k  
  
         t a s k   d a t a _ r e a d ( ) ;  
  
                 $ d i s p l a y ( " S c o r e b o a r d   r e a d " ) ;  
  
                 d r v 2 s b . g e t ( t x 1 ) ;  
                 m a i l 2 s b . g e t ( t x 2 ) ;  
  
                 t e m p _ a d d r   =   t x 1 . H a d d r [ 1 9 : 0 ] ;  
  
                 $ d i s p l a y ( " T e m p   a d d r e s s   =   % h " ,   t e m p _ a d d r ) ;  
                 $ d i s p l a y ( " R e a d   d a t a   f r o m   D U T   % h " ,   t x 2 . P r d a t a ) ;   / /   d a t a   f r o m   m o n i t o r / D U T  
                 $ d i s p l a y ( " D a t a   f r o m   T B   m e m o r y   % h " ,   m e m _ t b [ t e m p _ a d d r ] ) ;  
  
                 / /   A s s e r t   t h a t   t h e   d a t a   r e a d   m a t c h e s   t h e   d a t a   i n   t h e   m e m o r y   m o d e l  
                         a s s e r t   ( t x 2 . P r d a t a   = =   m e m _ t b [ t e m p _ a d d r ] )  
                         e l s e   $ e r r o r ( " D a t a   r e a d i n g   f a i l e d " ) ;  
  
                 $ d i s p l a y ( " " ) ;  
 	 # 1 0 ;  
         e n d t a s k  
  
 e n d c l a s s  
  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     T e s t  
 / /   F i l e :         t e s t . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 7 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   T e s t   c l a s s   f o r m s   t h e   b a c k b o n e   o f   a n y   t e s t b e n c h   i n   a   S y s t e m V e r i l o g    
 / /   v e r i f i c a t i o n   e n v i r o n m e n t .   T h i s   c l a s s   i n t e g r a t e s   a l l   t h e   t e s t   c a s e s   d e f i n e d    
 / /   i n   t h e   e n v i r o n m e n t   a n d   o r c h e s t r a t e s   t h e i r   e x e c u t i o n   o v e r   t h e   c o u r s e   o f   a    
 / /   s i m u l a t i o n   r u n .  
 / /  
 / /   I n   t h i s   p a r t i c u l a r   s c e n a r i o ,   t h e   T e s t   c l a s s   c r e a t e s   a n   i n s t a n c e   o f   t h e    
 / /   e n v i r o n m e n t   c l a s s ,   p r o v i d i n g   i t   w i t h   t h e   h a n d l e   t o   t h e   i n t e r f a c e   o b j e c t .    
 / /   T h e   ' r u n '   t a s k   o f   t h i s   c l a s s   s t a r t s   t h e   e n v i r o n m e n t   a n d   p e r f o r m s   t h e   t e s t    
 / /   s e q u e n c e s   r e p e a t e d l y   o v e r   m u l t i p l e   c l o c k   c y c l e s .    
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
 c l a s s   t e s t ;  
     e n v i r o n m e n t   e n v ;     / /   c r e a t e s   h a n d l e  
  
     f u n c t i o n   n e w ( v i r t u a l   a h b _ a p b _ b f m _ i f   i ) ;  
         e n v   =   n e w ( i ) ;    
     e n d f u n c t i o n   :   n e w  
      
     t a s k   r u n ( ) ;  
          
         $ d i s p l a y ( " i n   t e s t " ) ;        
         e n v . c r e a t e ( ) ;      
  
         r e p e a t ( 5 0 )                  
         b e g i n    
              
             $ d i s p l a y ( " i n   t e s t   r e p e a t " ) ;  
  
             e n v . e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 8 _ b y t e _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ w r a p 8 _ h a l f w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 8 _ w o r d _ n o n s e q _ w r a p 8 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 8 _ b y t e _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r 8 _ h a l f w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 8 _ w o r d _ n o n s e q _ i n c r 8 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ s i n g l e _ w o r d _ s e q _ s i n g l e _ H t r a n s f e r _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ s i n g l e _ b y t e _ s e q _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r _ h a l f w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r _ w o r d _ s e q _ i n c r _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 4 _ b y t e _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 4 _ w o r d _ s e q _ w r a p 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ b y t e _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ w o r d _ s e q _ i n c r 4 _ H b u r s t _ o k a y ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ s i n g l e _ b y t e _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ s i n g l e _ h a l f w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ s i n g l e _ w o r d _ n o n s e q _ s i n g l e _ H t r a n s f e r _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r _ b y t e _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r _ h a l f w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r _ w o r d _ n o n s e q _ i n c r _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 4 _ b y t e _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ w r a p 4 _ h a l f w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ w r a p 4 _ w o r d _ n o n s e q _ w r a p 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ b y t e _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ r e a d _ i n c r 4 _ h a l f w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ w o r d _ n o n s e q _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ w o r d _ i d l e _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ i n c r 4 _ w o r d _ b u s y _ i n c r 4 _ H b u r s t _ r e s e t ( ) ;  
             # 5 ;  
             e n v . e n v _ w r i t e _ s i n g l e _ b y t e _ i d l e _ s i n g l e _ H t r a n s f e r _ e r r o r ( ) ;  
             # 5 ;  
          
         e n d  
     e n d t a s k  
 e n d c l a s s  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     T o p - l e v e l   M o d u l e  
 / /   F i l e :         t o p . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 8 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   t o p - l e v e l   m o d u l e   o f   t h e   t e s t b e n c h ,   a h b _ a p b _ t o p ,   i n t e g r a t e s   a l l   t h e    
 / /   c o m p o n e n t s   o f   t h e   t e s t b e n c h   a n d   c o n n e c t s   t h e m   w i t h   t h e   D U T   ( D e v i c e   U n d e r    
 / /   V e r i f i c a t i o n ) .   T h e   D U T   i s   a n   A H B   t o   A P B   b r i d g e ,   a n d   i t s   m o d u l e   n a m e   i s    
 / /   ' B r i d g e _ T o p ' .  
 / /  
 / /   T h e   t o p   m o d u l e   i n c l u d e s   s e v e r a l   f i l e s :  
 / /   1 .   t r a n s a c t i o n s . s v   -   d e f i n e s   t h e   t r a n s a c t i o n   c l a s s  
 / /   2 .   g e n e r a t o r . s v   -   d e f i n e s   t h e   g e n e r a t o r   c l a s s  
 / /   3 .   i n t e r f a c e . s v   -   d e f i n e s   t h e   i n t e r f a c e   c l a s s  
 / /   4 .   d r i v e r . s v   -   d e f i n e s   t h e   d r i v e r   c l a s s  
 / /   5 .   m o n i t o r . s v   -   d e f i n e s   t h e   m o n i t o r   c l a s s  
 / /   6 .   s c o r e b o a r d . s v   -   d e f i n e s   t h e   s c o r e b o a r d   c l a s s  
 / /   7 .   c o v e r a g e . s v   -   d e f i n e s   t h e   c o v e r a g e   c o l l e c t o r   c l a s s  
 / /   8 .   e n v i r o n m e n t . s v   -   d e f i n e s   t h e   e n v i r o n m e n t   c l a s s  
 / /   9 .   t e s t . s v   -   d e f i n e s   t h e   t e s t   c l a s s  
 / /   1 0 .   b r i d g e _ t o p . v   -   t h i s   i s   p r e s u m a b l y   t h e   V e r i l o g   s o u r c e   c o d e   f o r   t h e   D U T  
 / /  
 / /   T h e   t o p   m o d u l e   a l s o   g e n e r a t e s   a   c l o c k   s i g n a l   ' c l k '   w i t h   a   p e r i o d   o f   1 0   n s    
 / /   ( h a l f   p e r i o d   o f   5   n s ) .   T h e   r e s e t   s i g n a l   ' r e s e t '   i s   i n i t i a l i z e d   t o   0   a n d   t h e n    
 / /   s e t   t o   1   a f t e r   1 0   t i m e   u n i t s .  
 / /  
 / /   T h e   t e s t   c l a s s   i s   i n s t a n t i a t e d   a s   ' t e s t _ h ' .   T h e   r u n   m e t h o d   o f   t h e   t e s t    
 / /   c l a s s   i s   c a l l e d   t o   s t a r t   t h e   t e s t .  
 / /  
 / /   T h e   s i m u l a t i o n   i s   s t o p p e d   a f t e r   1 0 0 0 0 0   t i m e   u n i t s   u s i n g   t h e   ' $ s t o p '    
 / /   s y s t e m   t a s k .  
 / /  
 / /   T h e   D U T   i s   i n s t a n t i a t e d   a s   ' d u t '   a n d   c o n n e c t e d   t o   t h e   t e s t b e n c h   u s i n g   a n    
 / /   i n s t a n c e   o f   t h e   a h b _ a p b _ b f m _ i f   i n t e r f a c e   n a m e d   ' b f m ' .   T h i s   i n t e r f a c e    
 / /   i n s t a n c e   i s   u s e d   t o   d r i v e   s i g n a l s   i n t o   t h e   D U T   a n d   m o n i t o r   s i g n a l s   c o m i n g    
 / /   f r o m   t h e   D U T .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
  
 ` i n c l u d e   " t r a n s a c t i o n s . s v "  
 ` i n c l u d e   " g e n e r a t o r . s v "  
 ` i n c l u d e   " i n t e r f a c e . s v "  
 ` i n c l u d e   " d r i v e r . s v "  
 ` i n c l u d e   " m o n i t o r . s v "  
 ` i n c l u d e   " s c o r e b o a r d . s v "  
 ` i n c l u d e   " c o v e r a g e . s v "  
 ` i n c l u d e   " e n v i r o n m e n t . s v "  
 ` i n c l u d e   " t e s t . s v "      
 ` i n c l u d e   " b r i d g e _ t o p . v "      
  
 m o d u l e   a h b _ a p b _ t o p ;  
  
     l o g i c   c l k ,   r e s e t ;  
  
     / /   G e n e r a t e s   c l k   w i t h   a   t i m e   p e r i o d   o f   5   n s  
     a l w a y s  
     b e g i n  
         f o r e v e r   b e g i n  
             # 5   c l k   =   ~ c l k ;  
         e n d  
     e n d  
  
    
  
     a h b _ a p b _ b f m _ i f   b f m ( c l k ,   r e s e t ) ;   / /   C o n n e c t   c l o c k   a n d   r e s e t  
  
  
     / /   C o n n e c t i n g   D U T   s i g n a l s   w i t h   s i g n a l s   p r e s e n t   o n   t h e   i n t e r f a c e  
 / /   C o n n e c t i n g   D U T   s i g n a l s   w i t h   s i g n a l s   p r e s e n t   o n   t h e   i n t e r f a c e  
 B r i d g e _ T o p   d u t (  
         . H c l k ( b f m . c l k ) ,  
         . H r e s e t n ( b f m . r e s e t n ) ,  
         . H w r i t e ( b f m . H w r i t e ) ,  
         . H r e a d y i n ( b f m . H r e a d y i n ) ,  
         . H t r a n s ( b f m . H t r a n s ) ,  
         . H w d a t a ( b f m . H w d a t a ) ,  
         . H a d d r ( b f m . H a d d r ) ,  
         . H r d a t a ( b f m . H r d a t a ) ,  
         . H r e s p ( b f m . H r e s p ) ,  
         . H r e a d y o u t ( b f m . H r e a d y o u t ) ,  
         . P r d a t a ( b f m . P r d a t a ) ,  
         . P w d a t a ( b f m . P w d a t a ) ,  
         . P a d d r ( b f m . P a d d r ) ,  
         . P s e l x ( b f m . P s e l x ) ,  
         . P w r i t e ( b f m . P w r i t e ) ,  
         . P e n a b l e ( b f m . P e n a b l e )  
 ) ;  
  
  
     / /   t e s t   a h b _ a p b _ t e s t ( b f m ) ;   / /   - >   n o t   i n i t i a l i z e d  
         t e s t   t e s t _ h ;  
         T r a n s a c t i o n   t r a n s ;  
     i n i t i a l   b e g i n  
         $ d i s p l a y ( " i n   t o p " ) ;  
         t r a n s   =   n e w ( ) ;  
         t r a n s . c o v _ c g . s a m p l e ( ) ;     / /   - >   t o   g e t   t h e   c o v e r a g e  
 	 t e s t _ h   =   n e w ( b f m ) ;  
 	 t e s t _ h . r u n ( ) ;  
  
 	  
     e n d  
  
   / /   I n i t i a l i z e   c l k   a n d   r e s e t  
     i n i t i a l   b e g i n  
         c l k   =   1 ;  
         r e s e t   =   0 ;  
         # 1 0  
         r e s e t   =   1 ;  
 	  
  
         # 1 0 0 0 0 0 ;  
         $ s t o p ;   / /   S t o p s   s i m u l a t i o n  
     e n d  
  
 e n d m o d u l e  
  
  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   P r o j e c t :   A H B   A P B   B r i d g e   V e r i f i c a t i o n  
 / /   M o d u l e :     T r a n s a c t i o n  
 / /   F i l e :         t r a n s a c t i o n s . s v  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 / /   A u t h o r :     M o h a m e d   G h o n i m  
 / /   C r e a t e d :   2 5 - J u l - 2 0 2 3  
 / /  
 / /   D e s c r i p t i o n :    
 / /   T h e   T r a n s a c t i o n   c l a s s   d e f i n e s   t h e   c h a r a c t e r i s t i c s   a n d   b e h a v i o r   o f   a    
 / /   t r a n s a c t i o n   t h a t   c a n   o c c u r   i n   t h e   A H B   A P B   B r i d g e .   E a c h   t r a n s a c t i o n   c o n t a i n s    
 / /   d e t a i l s   s u c h   a s   t h e   a d d r e s s ,   d a t a ,   t r a n s a c t i o n   t y p e ,   a n d   o t h e r   p r o p e r t i e s    
 / /   r e q u i r e d   f o r   A H B   a n d   A P B   p r o t o c o l s .   A   s e t   o f   c o n s t r a i n t s   i s   d e f i n e d   t o    
 / /   e n s u r e   v a l i d   t r a n s a c t i o n s   a r e   g e n e r a t e d .  
 / /    
 / /   T h i s   c l a s s   a l s o   f e a t u r e s   m e t h o d s   t o   u p d a t e   t r a n s a c t i o n   t y p e   b a s e d   o n   w h e t h e r    
 / /   a   r e a d   o r   w r i t e   o p e r a t i o n   i s   p e r f o r m e d ,   p r i n t   t h e   d e t a i l s   o f   t h e   t r a n s a c t i o n ,    
 / /   a n d   d e f i n e   a   c o v e r g r o u p   f o r   c o v e r a g e   c o l l e c t i o n .   T h e   c o v e r a g e   i s   m e a s u r e d    
 / /   f o r   v a r i o u s   o p e r a t i o n s ,   s i z e s ,   a n d   b u r s t   t y p e s   w h i c h   e n s u r e s   c o m p r e h e n s i v e    
 / /   v e r i f i c a t i o n .  
 / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
  
  
 c l a s s   T r a n s a c t i o n ;  
  
     t y p e d e f   e n u m   { A H B _ R E A D ,   A H B _ W R I T E }   t r a n s _ t y p e _ e ;  
     t r a n s _ t y p e _ e   t r a n s _ t y p e ;  
  
     r a n d c   b i t   [ 3 1 : 0 ]   H a d d r ;  
     r a n d c   b i t   [ 3 1 : 0 ]   H w d a t a ;  
     r a n d c   b i t   H w r i t e ;  
     r a n d c   b i t   [ 1 : 0 ]   H t r a n s ;  
     r a n d c   b i t   [ 2 : 0 ]   H s i z e ;  
     r a n d c   b i t   [ 2 : 0 ]   H b u r s t ;  
     r a n d c   b i t   [ 3 1 : 0 ]   P a d d r ;  
     r a n d c   b i t   [ 3 1 : 0 ]   P w d a t a ;  
     r a n d c   b i t   P w r i t e ;  
     r a n d c   b i t   [ 2 : 0 ]   P s e l x ;  
     r a n d c   b i t   h r e s p ; 	 / /   m a y   r e m o v e   l a t e r  
     r a n d c   b i t   h r e s e t ;     / /   R e s e t   s i g n a l  
  
     r a n d c   b i t   P e n a b l e ;     / /   A d d e d   t h i s   l i n e  
     r a n d c   b i t   [ 3 1 : 0 ]   P r d a t a ;   / / a d d e d   t h i s  
  
  
  
     c o n s t r a i n t   a d d r e s s   {  
         H a d d r [ 3 1 : 1 2 ]   = =   ' b 0 ;  
     }  
     c o n s t r a i n t   s i z e _ d a t a   { H s i z e   i n s i d e   { 0 , 1 , 2 } ; }  
     c o n s t r a i n t   b u r s t _ d a t a   { H b u r s t   i n s i d e   { 0 , 1 , 2 } ; }  
  
 c o v e r g r o u p   c o v _ c g ;       / /   - >   n o   @ ( H t r a n s . . . )   n o t   e v e n t s  
   	       H w r i t e _ c p :   c o v e r p o i n t   H w r i t e   {  
             	     b i n s   r e a d     =   { 1 ' b 0 } ;  
             	     b i n s   w r i t e   =   { 1 ' b 1 } ;  
                 }  
                 H t r a n s _ c p :   c o v e r p o i n t   H t r a n s   {  
                         b i n s   n o n _ s e q   =   { 2 ' b 1 0 } ;  
                         b i n s   i d l e         =   { 2 ' b 0 0 } ;  
                         b i n s   s e q           =   { 2 ' b 1 1 } ;  
                         / / b i n s   b u s y         =   { 2 ' b 0 1 } ;  
                 }  
                 H s i z e _ c p :   c o v e r p o i n t   H s i z e   {  
                         b i n s   s i z e _ b y t e           =   { 3 ' b 0 0 0 } ;  
                         b i n s   s i z e _ h a l f w o r d   =   { 3 ' b 0 0 1 } ;  
                         b i n s   s i z e _ w o r d           =   { 3 ' b 0 1 0 } ;  
                 }  
                 H b u r s t _ c p :   c o v e r p o i n t   H b u r s t   {  
                         b i n s   s i n g l e   =   { 3 ' b 0 0 0 } ;  
                         b i n s   i n c r       =   { 3 ' b 0 0 1 } ;  
                         b i n s   w r a p 4     =   { 3 ' b 0 1 0 } ;  
                         b i n s   i n c r 4     =   { 3 ' b 0 1 1 } ;  
                 }  
                 / /   C r o s s   c o v e r a g e  
         H w r i t e _ x _ h t r a n s :   c r o s s   H w r i t e _ c p ,   H t r a n s _ c p ;  
         H w r i t e _ x _ h s i z e :   c r o s s   H w r i t e _ c p ,   H s i z e _ c p ;  
         H w r i t e _ x _ h b u r s t :   c r o s s   H w r i t e _ c p ,   H b u r s t _ c p ;  
         e n d g r o u p  
  
     f u n c t i o n   n e w ( ) ;  
         c o v _ c g   =   n e w ;  
     e n d f u n c t i o n  
  
     f u n c t i o n   v o i d   u p d a t e _ t r a n s _ t y p e ( ) ;  
         i f   ( H w r i t e   = =   1 )    
             t r a n s _ t y p e   =   T r a n s a c t i o n : : A H B _ W R I T E ;  
         e l s e  
             t r a n s _ t y p e   =   T r a n s a c t i o n : : A H B _ R E A D ;  
  
         / /   C a l l   c o v _ c g . s a m p l e ( )   h e r e   a f t e r   t h e   t r a n s _ t y p e   i s   u p d a t e d  
         c o v _ c g . s a m p l e ( ) ;  
     e n d f u n c t i o n  
  
     f u n c t i o n   v o i d   p r i n t _ t r a n s a c t i o n ( ) ;  
         $ d i s p l a y ( " T r a n s a c t i o n   D e t a i l s : " ) ;  
         $ d i s p l a y ( " - - - - - - - - - - - - - - - - - - - " ) ;  
         $ d i s p l a y ( " T r a n s a c t i o n   T y p e :   % s " ,   t r a n s _ t y p e . n a m e ( ) ) ;  
         $ d i s p l a y ( " H a d d r :   % 0 d " ,   H a d d r ) ;  
         $ d i s p l a y ( " H w d a t a :   % 0 d " ,   H w d a t a ) ;  
         $ d i s p l a y ( " H w r i t e :   % 0 b " ,   H w r i t e ) ;  
         $ d i s p l a y ( " H t r a n s :   % 0 b " ,   H t r a n s ) ;  
         $ d i s p l a y ( " H s i z e :   % 0 b " ,   H s i z e ) ;  
         $ d i s p l a y ( " H b u r s t :   % 0 b " ,   H b u r s t ) ;  
         $ d i s p l a y ( " P a d d r :   % 0 d " ,   P a d d r ) ;  
         $ d i s p l a y ( " P w d a t a :   % 0 d " ,   P w d a t a ) ;  
         $ d i s p l a y ( " P w r i t e :   % 0 b " ,   P w r i t e ) ;  
         $ d i s p l a y ( " P s e l x :   % 0 b " ,   P s e l x ) ;  
         $ d i s p l a y ( " P e n a b l e :   % 0 b " ,   P e n a b l e ) ;  
     e n d f u n c t i o n  
  
      
  
 e n d c l a s s  
 